** Profile: "Startup_TB-trans"  [ c:\elab_model_ws\elab_model_ds\part_numbers\tps61322\release_ti\pspice\tps61322_pspice_trans\tps61322_trans-pspicefiles\startup_tb\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tps61322_trans.lib" 
* From [PSPICE NETLIST] section of C:\Users\a0132703\Documents\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "C:\Cadence\SPB_166\tools\pspice\library\nom.lib" 

*Analysis directives: 
.TRAN  0 1.5m 0 10n SKIPBP 
.OPTIONS ADVCONV
.OPTIONS ITL2= 40
.OPTIONS ITL4= 40
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\Startup_TB.net" 


.END
